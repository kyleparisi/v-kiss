module main

fn hello() string {
	return "Hello, Testing!"
}

fn main() {
	println(hello())
}
